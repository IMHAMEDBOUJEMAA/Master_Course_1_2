library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UAL_4bits is
port( A, B: in std_logic_vector(3 downto 0);
      op: in std_logic_vector(2 downto 0);
      R: out std_logic_vector(3 downto 0));
end entity UAL_4bits;

architecture Behavioral of UAL_4bits is
begin
  process(A, B, op)
  begin
    case op is
      when "000" =>
        R <= std_logic_vector(unsigned(A) + unsigned(B));
      when "001" =>
        R <= std_logic_vector(unsigned(A) - unsigned(B));
      when "010" =>
        R <= std_logic_vector(unsigned(A) + 1);
      when "011" =>
        R <= std_logic_vector(unsigned(A) - 1);
      when "100" =>
        R <= A and B;
      when "101" =>
        R <= A or B;
      when "110" =>
        R <= not A;
      when "111" =>
        R <= A xor B;
      when others =>
        R <= (others => '0');
    end case;
  end process;
end architecture Behavioral;

