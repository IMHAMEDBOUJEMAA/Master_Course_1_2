-- 4 bit FULL ADDER
-- Entity 
entity FULLADD4 is 
port (a0, b0, a1, b1, a2, b2, a3, b3, c0 : in bit;
	c4, s0, s1,s2,s3 : out bit);
end FULLADD4;

--Architecture 
architecture struct of FULLADD4 is 
-- signals 
signal c1, c2, c3 : bit;
-- use 1 bit FULL ADDER
component FULLADD 
port (A,B,CIN : in bit ; S,COUT : out bit);
end component;
-- Begin 

begin
 
FA1:FULLADD port map (a0,b0,c0,s0,c1);
FA2:FULLADD port map (a1,b1,c1,s1,c2);
FA3:FULLADD port map (a2,b2,c2,s2,c3);
FA4:FULLADD port map (a3,b3,c3,s3,c4);
end struct; 